/*
 * cursor_uart_tx.v
 *
 * Instrument-Grade UART Transmitter for Boreal Neuro-Core.
 * Packet Frame (6 bytes):
 * [0] SYNC (0xAA)
 * [1] VERSION(2) | BUTTONS(2) | SAFETY(4)
 * [2] DX (signed 8-bit)
 * [3] DY (signed 8-bit)
 * [4] FRAME_ID (8-bit counter)
 * [5] CRC8 (Poly 0x07)
 */
module cursor_uart_tx #(
    parameter CLKS_PER_BIT = 217
)(
    input  wire        clk,
    input  wire        rst,
    input  wire        send,
    input  wire [1:0]  buttons,
    input  wire signed [7:0] dx,
    input  wire signed [7:0] dy,
    input  wire [7:0]  frame_id,
    input  wire [3:0]  safety_flags,
    output reg         tx,
    output reg         tx_busy
);

    localparam VERSION = 2'b01;

    reg [7:0]  packet [0:5];
    reg [2:0]  byte_idx;
    reg [3:0]  bit_idx;
    reg [15:0] clk_cnt;
    reg        sending;

    // CRC8 Calculation (Combinatorial for the frame)
    function [7:0] crc8;
        input [39:0] data; // 5 bytes
        integer i;
        reg [7:0] crc;
        begin
            crc = 8'h00;
            for (i = 39; i >= 0; i = i - 1) begin
                if ((crc[7] ^ data[i]) == 1'b1)
                    crc = (crc << 1) ^ 8'h07;
                else
                    crc = (crc << 1);
            end
            crc8 = crc;
        end
    endfunction

    wire [7:0] vbs = {VERSION, buttons, safety_flags};
    wire [7:0] final_crc = crc8({vbs, dx, dy, frame_id, 8'h00}); // Placeholder logic for demonstration

    // Simple XOR for now to ensure bitwise stability in the FSM before full expansion
    // Using blocking assignments for the checksum to avoid the race condition
    reg [7:0] checksum_calc;

    always @(posedge clk) begin
        if (rst) begin
            tx <= 1;
            sending <= 0;
            tx_busy <= 0;
            byte_idx <= 0;
            bit_idx <= 0;
            clk_cnt <= 0;
        end else if (send && !sending) begin
            packet[0] <= 8'hAA;
            packet[1] <= vbs;
            packet[2] <= dx;
            packet[3] <= dy;
            packet[4] <= frame_id;
            // Formal CRC8 calculation over bytes 1 to 4
            packet[5] <= crc8({vbs, dx, dy, frame_id, 8'h00}); 

            byte_idx <= 0;
            bit_idx <= 0;
            clk_cnt <= 0;
            sending <= 1;
            tx_busy <= 1;
        end else if (sending) begin
            if (clk_cnt == CLKS_PER_BIT - 1) begin
                clk_cnt <= 0;
                if (bit_idx == 0) begin
                    tx <= 0; // Start
                    bit_idx <= 1;
                end else if (bit_idx <= 8) begin
                    tx <= packet[byte_idx][bit_idx-1];
                    bit_idx <= bit_idx + 1;
                end else begin
                    tx <= 1; // Stop
                    bit_idx <= 0;
                    if (byte_idx == 5) begin
                        sending <= 0;
                        tx_busy <= 0;
                    end else begin
                        byte_idx <= byte_idx + 1;
                    end
                end
            end else begin
                clk_cnt <= clk_cnt + 1;
            end
        end
    end

endmodule
